library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity OPCODEM is
    Generic( 
        m : integer := 5;
        n : integer := 20
        );
    Port(
        OPCODE : in STD_LOGIC_VECTOR(m-1 downto 0);
        MIC : out STD_LOGIC_VECTOR(n-1 downto 0)
    );
end OPCODEM;

architecture A_OPCODEM of OPCODEM is

TYPE BANCO IS ARRAY (0 to (2**m)-1) of std_logic_vector(n-1 downto 0);       
CONSTANT DEFAULT_MOP : BANCO :=(
    "00000100000001110001", --Verificacion
    "00000000100000000000", --LI
    "00001000100000001000", --LWI
    "00000100000000001100", --SWI
    "00000100011000110101", --SW
    "00001000101000110011", --ADDI
    "00001000101001110011", --SUBI
    "00001000101000000011", --ANDI
    "00001000101000010011", --ORI
    "00001000101000100011", --XORI
    "00001000101011010011", --NANDI
    "00001000101011000011", --NORI
    "00001000101001100011", --XNORI
    "00110000001100110011", --BEQI
    "00110000001100110011", --BNEI
    "00110000001100110011", --BLTI
    "00110000001100110011", --BLETI
    "00110000001100110011", --BGTI
    "00110000001100110011", --BGETI
    "00100000000000000000", --B
    "10100000000000000000", --CALL
    "01100000000000000000", --RET
    "00000000000000000000", --NOP
    "00001000111000110001", --LW
    others => (others => '0')
    );
    
begin
    MIC <= DEFAULT_MOP(conv_integer(OPCODE));
end A_OPCODEM;
